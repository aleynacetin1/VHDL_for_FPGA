library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity and_component is
    Port ( a : in STD_LOGIC;
           b : in STD_LOGIC;
           c : out STD_LOGIC);
end and_component;

architecture Behavioral of and_component is

begin
    c <= a and b;

end Behavioral;
